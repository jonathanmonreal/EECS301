module speed_counter();

endmodule