module brake(clock, brake, l_signal, r_signal, l_lights, c_lights, r_lights);

endmodule