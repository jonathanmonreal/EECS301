module speed_counter(input_a, input_b, speed);

	input input_a, input_b;
	output speed;

endmodule