// Jonathan Monreal
// This module is a simple clock divider

module button_clock(clk, clk_out);

	input clk;
	output wire clk_out;
	
	reg [16:0] counter =17'b0;
	// The output is the msb of the counter
	assign clk_out = counter[16];
	
	always @(posedge clk)
		begin
			counter <= counter + 1'b1;
		end
		
endmodule