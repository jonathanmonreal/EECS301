module pwm();
endmodule